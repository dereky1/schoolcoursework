library IEEE;
use IEEE.STD_LOGIC_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity alu32 is
port(
	A : in std_logic_vector(31 downto 0);
	B : in std_logic_vector(31 downto 0);
	alu_op : in std_logic_vector(3 downto 0);
	g : out std_logic;
	e : out std_logic;
	l : out std_logic;
	output : out std_logic_vector(31 downto 0);
	cout : inout std_logic;
	over : out std_logic
);
end alu32;

architecture data of alu32 is
component alu_1bit IS
PORT (
A : IN STD_LOGIC ;
B : IN STD_LOGIC ;
cin : IN STD_LOGIC ;
alu_op : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
output : OUT STD_LOGIC ;
cout : OUT STD_LOGIC
);
END component alu_1bit ;

component carry_gen IS
PORT (
alu_op : IN std_logic_vector(3 downto 0) ;
cout : OUT std_logic
);
END component carry_gen ;

component comparator IS
PORT (
	in_0 : IN STD_LOGIC_vector (31 downto 0) ;
	in_1 : IN STD_LOGIC_vector (31 downto 0) ;
	greater : OUT STD_LOGIC ;
	equal : OUT STD_LOGIC ;
	less : OUT STD_LOGIC
);
END component comparator ;

signal c_intermediate : std_logic_vector(32 downto 0);
signal gc, ec, lc : std_logic;

begin

cm: comparator port map (A, B, gc, ec, lc);
cg: carry_gen port map (alu_op, c_intermediate(0));

alu_32_bit: for i in 0 to 31 generate

U0: alu_1bit port map (A(i),B(i),c_intermediate(i), alu_op, output(i), c_intermediate(i+1));

end generate alu_32_bit;

g <= '0' when alu_op <= "0100" else gc;
e <= '0' when alu_op <= "0100" else ec;
l <= '1' when alu_op <= "0100" else lc;

cout<= c_intermediate(32);	

over<= c_intermediate(31) xor c_intermediate(30); 

end data;